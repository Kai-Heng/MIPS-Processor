------------------------------------
-- Kai Heng Gan
-- Cyber Security Engineering
-- Iowa State University
------------------------------------

--decoder.vhd

library IEEE;
use IEEE.std_logic_1164.all;

entity decoder5to32 is
  port(WA	: in std_logic_vector(4 downto 0);
       En        : in std_logic;
       Q          : out std_logic_vector(31 downto 0));   -- Data value output   

end decoder5to32;

architecture dataflow of decoder5to32 is
begin

  process (WA)
    begin
	case WA is
		when "00000" => Q <= "00000000000000000000000000000001"; -- $0
		when "00001" => Q <= "00000000000000000000000000000010"; -- $1
		when "00010" => Q <= "00000000000000000000000000000100"; -- $2
		when "00011" => Q <= "00000000000000000000000000001000"; -- $3
		when "00100" => Q <= "00000000000000000000000000010000"; -- $4
		when "00101" => Q <= "00000000000000000000000000100000"; -- $5
		when "00110" => Q <= "00000000000000000000000001000000"; -- $6
		when "00111" => Q <= "00000000000000000000000010000000"; -- $7
		when "01000" => Q <= "00000000000000000000000100000000"; -- $8
		when "01001" => Q <= "00000000000000000000001000000000"; -- $9
		when "01010" => Q <= "00000000000000000000010000000000"; -- $10
		when "01011" => Q <= "00000000000000000000100000000000"; -- $11
		when "01100" => Q <= "00000000000000000001000000000000"; -- $12
		when "01101" => Q <= "00000000000000000010000000000000"; -- $13
		when "01110" => Q <= "00000000000000000100000000000000"; -- $14
		when "01111" => Q <= "00000000000000001000000000000000"; -- $15
		when "10000" => Q <= "00000000000000010000000000000000"; -- $16
		when "10001" => Q <= "00000000000000100000000000000000"; -- $17
		when "10010" => Q <= "00000000000001000000000000000000"; -- $18
		when "10011" => Q <= "00000000000010000000000000000000"; -- $19
		when "10100" => Q <= "00000000000100000000000000000000"; -- $20
		when "10101" => Q <= "00000000001000000000000000000000"; -- $21
		when "10110" => Q <= "00000000010000000000000000000000"; -- $22
		when "10111" => Q <= "00000000100000000000000000000000"; -- $23
		when "11000" => Q <= "00000001000000000000000000000000"; -- $24
		when "11001" => Q <= "00000010000000000000000000000000"; -- $25
		when "11010" => Q <= "00000100000000000000000000000000"; -- $26
		when "11011" => Q <= "00001000000000000000000000000000"; -- $27
		when "11100" => Q <= "00010000000000000000000000000000"; -- $28
		when "11101" => Q <= "00100000000000000000000000000000"; -- $29
		when "11110" => Q <= "01000000000000000000000000000000"; -- $30
		when "11111" => Q <= "10000000000000000000000000000000"; -- $31
		when others => Q <= "00000000000000000000000000000000";
	end case;
  end process;
  
end dataflow;